`timescale 1ns / 1ps



module two_bit_or(
        input A,B,
        output Y
    );
    assign Y = A|B;
endmodule
